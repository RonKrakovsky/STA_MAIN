/* 
RON KRAKOVSKY
out = log10(in) ufix(25,7) = 32*/

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--------------------------------------------------

entity Log_10 is
port(	
	csi_sink_clk	 	 : in std_logic; -- clock
	rsi_sink_reset	 	 : in std_logic; -- reset in LOW = '0'
	i_bit_index			 : in std_logic_vector(31 downto 0);
	o_bit_index			 : out std_logic_vector(31 downto 0);
	asi_sink_data		 : in std_logic_vector(30 downto 0); --ufix31_En3
	aso_source_data		 : out unsigned(31 downto 0) --ufix32_En7
);
end Log_10;  


--------------------------------------------------

architecture behav of Log_10 is
signal bit_fft_index : std_logic_vector(31 downto 0);
begin
	process(csi_sink_clk, rsi_sink_reset)
    begin
		if rsi_sink_reset = '0' then 
			aso_source_data <= (others => '0');
		elsif rising_edge(csi_sink_clk) then 
			bit_fft_index <= i_bit_index;
		
			case to_integer(unsigned(asi_sink_data)) is
when  0  to  8 => aso_source_data <= to_unsigned( 0 ,32);
when  9  to  9 => aso_source_data <= to_unsigned( 7 ,32);
when  10  to  10 => aso_source_data <= to_unsigned( 12 ,32);
when  11  to  11 => aso_source_data <= to_unsigned( 17 ,32);
when  12  to  12 => aso_source_data <= to_unsigned( 23 ,32);
when  13  to  13 => aso_source_data <= to_unsigned( 28 ,32);
when  14  to  14 => aso_source_data <= to_unsigned( 32 ,32);
when  15  to  15 => aso_source_data <= to_unsigned( 35 ,32);
when  16  to  16 => aso_source_data <= to_unsigned( 39 ,32);
when  17  to  17 => aso_source_data <= to_unsigned( 42 ,32);
when  18  to  18 => aso_source_data <= to_unsigned( 46 ,32);
when  19  to  19 => aso_source_data <= to_unsigned( 48 ,32);
when  20  to  20 => aso_source_data <= to_unsigned( 51 ,32);
when  21  to  21 => aso_source_data <= to_unsigned( 53 ,32);
when  22  to  22 => aso_source_data <= to_unsigned( 56 ,32);
when  23  to  23 => aso_source_data <= to_unsigned( 58 ,32);
when  24  to  24 => aso_source_data <= to_unsigned( 61 ,32);
when  25  to  25 => aso_source_data <= to_unsigned( 64 ,32);
when  26  to  27 => aso_source_data <= to_unsigned( 66 ,32);
when  28  to  29 => aso_source_data <= to_unsigned( 70 ,32);
when  30  to  31 => aso_source_data <= to_unsigned( 74 ,32);
when  32  to  33 => aso_source_data <= to_unsigned( 78 ,32);
when  34  to  34 => aso_source_data <= to_unsigned( 80 ,32);
when  35  to  36 => aso_source_data <= to_unsigned( 83 ,32);
when  37  to  38 => aso_source_data <= to_unsigned( 85 ,32);
when  39  to  40 => aso_source_data <= to_unsigned( 88 ,32);
when  41  to  41 => aso_source_data <= to_unsigned( 90 ,32);
when  42  to  43 => aso_source_data <= to_unsigned( 93 ,32);
when  44  to  46 => aso_source_data <= to_unsigned( 96 ,32);
when  47  to  48 => aso_source_data <= to_unsigned( 98 ,32);
when  49  to  50 => aso_source_data <= to_unsigned( 101 ,32);
when  51  to  52 => aso_source_data <= to_unsigned( 103 ,32);
when  53  to  55 => aso_source_data <= to_unsigned( 106 ,32);
when  56  to  57 => aso_source_data <= to_unsigned( 108 ,32);
when  58  to  60 => aso_source_data <= to_unsigned( 111 ,32);
when  61  to  63 => aso_source_data <= to_unsigned( 113 ,32);
when  64  to  66 => aso_source_data <= to_unsigned( 116 ,32);
when  67  to  69 => aso_source_data <= to_unsigned( 119 ,32);
when  70  to  72 => aso_source_data <= to_unsigned( 121 ,32);
when  73  to  76 => aso_source_data <= to_unsigned( 124 ,32);
when  77  to  80 => aso_source_data <= to_unsigned( 126 ,32);
when  81  to  83 => aso_source_data <= to_unsigned( 129 ,32);
when  84  to  87 => aso_source_data <= to_unsigned( 131 ,32);
when  88  to  91 => aso_source_data <= to_unsigned( 134 ,32);
when  92  to  96 => aso_source_data <= to_unsigned( 136 ,32);
when  97  to  100 => aso_source_data <= to_unsigned( 139 ,32);
when  101  to  105 => aso_source_data <= to_unsigned( 142 ,32);
when  106  to  110 => aso_source_data <= to_unsigned( 144 ,32);
when  111  to  115 => aso_source_data <= to_unsigned( 147 ,32);
when  116  to  121 => aso_source_data <= to_unsigned( 149 ,32);
when  122  to  126 => aso_source_data <= to_unsigned( 152 ,32);
when  127  to  132 => aso_source_data <= to_unsigned( 154 ,32);
when  133  to  139 => aso_source_data <= to_unsigned( 157 ,32);
when  140  to  145 => aso_source_data <= to_unsigned( 160 ,32);
when  146  to  152 => aso_source_data <= to_unsigned( 162 ,32);
when  153  to  159 => aso_source_data <= to_unsigned( 165 ,32);
when  160  to  167 => aso_source_data <= to_unsigned( 167 ,32);
when  168  to  175 => aso_source_data <= to_unsigned( 170 ,32);
when  176  to  183 => aso_source_data <= to_unsigned( 172 ,32);
when  184  to  191 => aso_source_data <= to_unsigned( 175 ,32);
when  192  to  200 => aso_source_data <= to_unsigned( 177 ,32);
when  201  to  210 => aso_source_data <= to_unsigned( 180 ,32);
when  211  to  220 => aso_source_data <= to_unsigned( 183 ,32);
when  221  to  230 => aso_source_data <= to_unsigned( 185 ,32);
when  231  to  241 => aso_source_data <= to_unsigned( 188 ,32);
when  242  to  252 => aso_source_data <= to_unsigned( 190 ,32);
when  253  to  264 => aso_source_data <= to_unsigned( 193 ,32);
when  265  to  277 => aso_source_data <= to_unsigned( 195 ,32);
when  278  to  290 => aso_source_data <= to_unsigned( 198 ,32);
when  291  to  304 => aso_source_data <= to_unsigned( 200 ,32);
when  305  to  318 => aso_source_data <= to_unsigned( 203 ,32);
when  319  to  333 => aso_source_data <= to_unsigned( 206 ,32);
when  334  to  349 => aso_source_data <= to_unsigned( 208 ,32);
when  350  to  365 => aso_source_data <= to_unsigned( 211 ,32);
when  366  to  382 => aso_source_data <= to_unsigned( 213 ,32);
when  383  to  400 => aso_source_data <= to_unsigned( 216 ,32);
when  401  to  419 => aso_source_data <= to_unsigned( 218 ,32);
when  420  to  439 => aso_source_data <= to_unsigned( 221 ,32);
when  440  to  460 => aso_source_data <= to_unsigned( 224 ,32);
when  461  to  482 => aso_source_data <= to_unsigned( 226 ,32);
when  483  to  504 => aso_source_data <= to_unsigned( 229 ,32);
when  505  to  528 => aso_source_data <= to_unsigned( 231 ,32);
when  529  to  553 => aso_source_data <= to_unsigned( 234 ,32);
when  554  to  579 => aso_source_data <= to_unsigned( 236 ,32);
when  580  to  606 => aso_source_data <= to_unsigned( 239 ,32);
when  607  to  635 => aso_source_data <= to_unsigned( 241 ,32);
when  636  to  665 => aso_source_data <= to_unsigned( 244 ,32);
when  666  to  696 => aso_source_data <= to_unsigned( 247 ,32);
when  697  to  729 => aso_source_data <= to_unsigned( 249 ,32);
when  730  to  763 => aso_source_data <= to_unsigned( 252 ,32);
when  764  to  800 => aso_source_data <= to_unsigned( 254 ,32);
when  801  to  837 => aso_source_data <= to_unsigned( 257 ,32);
when  838  to  877 => aso_source_data <= to_unsigned( 259 ,32);
when  878  to  918 => aso_source_data <= to_unsigned( 262 ,32);
when  919  to  961 => aso_source_data <= to_unsigned( 264 ,32);
when  962  to  1007 => aso_source_data <= to_unsigned( 267 ,32);
when  1008  to  1054 => aso_source_data <= to_unsigned( 270 ,32);
when  1055  to  1104 => aso_source_data <= to_unsigned( 272 ,32);
when  1105  to  1156 => aso_source_data <= to_unsigned( 275 ,32);
when  1157  to  1210 => aso_source_data <= to_unsigned( 277 ,32);
when  1211  to  1267 => aso_source_data <= to_unsigned( 280 ,32);
when  1268  to  1327 => aso_source_data <= to_unsigned( 282 ,32);
when  1328  to  1390 => aso_source_data <= to_unsigned( 285 ,32);
when  1391  to  1455 => aso_source_data <= to_unsigned( 287 ,32);
when  1456  to  1524 => aso_source_data <= to_unsigned( 290 ,32);
when  1525  to  1596 => aso_source_data <= to_unsigned( 293 ,32);
when  1597  to  1671 => aso_source_data <= to_unsigned( 295 ,32);
when  1672  to  1750 => aso_source_data <= to_unsigned( 298 ,32);
when  1751  to  1832 => aso_source_data <= to_unsigned( 300 ,32);
when  1833  to  1919 => aso_source_data <= to_unsigned( 303 ,32);
when  1920  to  2009 => aso_source_data <= to_unsigned( 305 ,32);
when  2010  to  2104 => aso_source_data <= to_unsigned( 308 ,32);
when  2105  to  2203 => aso_source_data <= to_unsigned( 311 ,32);
when  2204  to  2307 => aso_source_data <= to_unsigned( 313 ,32);
when  2308  to  2415 => aso_source_data <= to_unsigned( 316 ,32);
when  2416  to  2529 => aso_source_data <= to_unsigned( 318 ,32);
when  2530  to  2649 => aso_source_data <= to_unsigned( 321 ,32);
when  2650  to  2773 => aso_source_data <= to_unsigned( 323 ,32);
when  2774  to  2904 => aso_source_data <= to_unsigned( 326 ,32);
when  2905  to  3041 => aso_source_data <= to_unsigned( 328 ,32);
when  3042  to  3184 => aso_source_data <= to_unsigned( 331 ,32);
when  3185  to  3334 => aso_source_data <= to_unsigned( 334 ,32);
when  3335  to  3492 => aso_source_data <= to_unsigned( 336 ,32);
when  3493  to  3656 => aso_source_data <= to_unsigned( 339 ,32);
when  3657  to  3829 => aso_source_data <= to_unsigned( 341 ,32);
when  3830  to  4009 => aso_source_data <= to_unsigned( 344 ,32);
when  4010  to  4198 => aso_source_data <= to_unsigned( 346 ,32);
when  4199  to  4396 => aso_source_data <= to_unsigned( 349 ,32);
when  4397  to  4603 => aso_source_data <= to_unsigned( 351 ,32);
when  4604  to  4820 => aso_source_data <= to_unsigned( 354 ,32);
when  4821  to  5047 => aso_source_data <= to_unsigned( 357 ,32);
when  5048  to  5285 => aso_source_data <= to_unsigned( 359 ,32);
when  5286  to  5534 => aso_source_data <= to_unsigned( 362 ,32);
when  5535  to  5795 => aso_source_data <= to_unsigned( 364 ,32);
when  5796  to  6068 => aso_source_data <= to_unsigned( 367 ,32);
when  6069  to  6354 => aso_source_data <= to_unsigned( 369 ,32);
when  6355  to  6654 => aso_source_data <= to_unsigned( 372 ,32);
when  6655  to  6967 => aso_source_data <= to_unsigned( 375 ,32);
when  6968  to  7296 => aso_source_data <= to_unsigned( 377 ,32);
when  7297  to  7639 => aso_source_data <= to_unsigned( 380 ,32);
when  7640  to  7999 => aso_source_data <= to_unsigned( 382 ,32);
when  8000  to  8377 => aso_source_data <= to_unsigned( 385 ,32);
when  8378  to  8771 => aso_source_data <= to_unsigned( 387 ,32);
when  8772  to  9185 => aso_source_data <= to_unsigned( 390 ,32);
when  9186  to  9618 => aso_source_data <= to_unsigned( 392 ,32);
when  9619  to  10071 => aso_source_data <= to_unsigned( 395 ,32);
when  10072  to  10546 => aso_source_data <= to_unsigned( 398 ,32);
when  10547  to  11043 => aso_source_data <= to_unsigned( 400 ,32);
when  11044  to  11563 => aso_source_data <= to_unsigned( 403 ,32);
when  11564  to  12108 => aso_source_data <= to_unsigned( 405 ,32);
when  12109  to  12679 => aso_source_data <= to_unsigned( 408 ,32);
when  12680  to  13276 => aso_source_data <= to_unsigned( 410 ,32);
when  13277  to  13902 => aso_source_data <= to_unsigned( 413 ,32);
when  13903  to  14557 => aso_source_data <= to_unsigned( 415 ,32);
when  14558  to  15243 => aso_source_data <= to_unsigned( 418 ,32);
when  15244  to  15962 => aso_source_data <= to_unsigned( 421 ,32);
when  15963  to  16714 => aso_source_data <= to_unsigned( 423 ,32);
when  16715  to  17502 => aso_source_data <= to_unsigned( 426 ,32);
when  17503  to  18326 => aso_source_data <= to_unsigned( 428 ,32);
when  18327  to  19190 => aso_source_data <= to_unsigned( 431 ,32);
when  19191  to  20095 => aso_source_data <= to_unsigned( 433 ,32);
when  20096  to  21042 => aso_source_data <= to_unsigned( 436 ,32);
when  21043  to  22033 => aso_source_data <= to_unsigned( 439 ,32);
when  22034  to  23072 => aso_source_data <= to_unsigned( 441 ,32);
when  23073  to  24159 => aso_source_data <= to_unsigned( 444 ,32);
when  24160  to  25298 => aso_source_data <= to_unsigned( 446 ,32);
when  25299  to  26490 => aso_source_data <= to_unsigned( 449 ,32);
when  26491  to  27738 => aso_source_data <= to_unsigned( 451 ,32);
when  27739  to  29046 => aso_source_data <= to_unsigned( 454 ,32);
when  29047  to  30415 => aso_source_data <= to_unsigned( 456 ,32);
when  30416  to  31848 => aso_source_data <= to_unsigned( 459 ,32);
when  31849  to  33349 => aso_source_data <= to_unsigned( 462 ,32);
when  33350  to  34921 => aso_source_data <= to_unsigned( 464 ,32);
when  34922  to  36567 => aso_source_data <= to_unsigned( 467 ,32);
when  36568  to  38290 => aso_source_data <= to_unsigned( 469 ,32);
when  38291  to  40094 => aso_source_data <= to_unsigned( 472 ,32);
when  40095  to  41984 => aso_source_data <= to_unsigned( 474 ,32);
when  41985  to  43963 => aso_source_data <= to_unsigned( 477 ,32);
when  43964  to  46035 => aso_source_data <= to_unsigned( 479 ,32);
when  46036  to  48204 => aso_source_data <= to_unsigned( 482 ,32);
when  48205  to  50476 => aso_source_data <= to_unsigned( 485 ,32);
when  50477  to  52855 => aso_source_data <= to_unsigned( 487 ,32);
when  52856  to  55346 => aso_source_data <= to_unsigned( 490 ,32);
when  55347  to  57954 => aso_source_data <= to_unsigned( 492 ,32);
when  57955  to  60686 => aso_source_data <= to_unsigned( 495 ,32);
when  60687  to  63546 => aso_source_data <= to_unsigned( 497 ,32);
when  63547  to  66541 => aso_source_data <= to_unsigned( 500 ,32);
when  66542  to  69677 => aso_source_data <= to_unsigned( 503 ,32);
when  69678  to  72960 => aso_source_data <= to_unsigned( 505 ,32);
when  72961  to  76399 => aso_source_data <= to_unsigned( 508 ,32);
when  76400  to  79999 => aso_source_data <= to_unsigned( 510 ,32);
when  80000  to  83770 => aso_source_data <= to_unsigned( 513 ,32);
when  83771  to  87718 => aso_source_data <= to_unsigned( 515 ,32);
when  87719  to  91852 => aso_source_data <= to_unsigned( 518 ,32);
when  91853  to  96181 => aso_source_data <= to_unsigned( 520 ,32);
when  96182  to  100714 => aso_source_data <= to_unsigned( 523 ,32);
when  100715  to  105460 => aso_source_data <= to_unsigned( 526 ,32);
when  105461  to  110430 => aso_source_data <= to_unsigned( 528 ,32);
when  110431  to  115635 => aso_source_data <= to_unsigned( 531 ,32);
when  115636  to  121084 => aso_source_data <= to_unsigned( 533 ,32);
when  121085  to  126791 => aso_source_data <= to_unsigned( 536 ,32);
when  126792  to  132766 => aso_source_data <= to_unsigned( 538 ,32);
when  132767  to  139024 => aso_source_data <= to_unsigned( 541 ,32);
when  139025  to  145576 => aso_source_data <= to_unsigned( 543 ,32);
when  145577  to  152436 => aso_source_data <= to_unsigned( 546 ,32);
when  152437  to  159620 => aso_source_data <= to_unsigned( 549 ,32);
when  159621  to  167143 => aso_source_data <= to_unsigned( 551 ,32);
when  167144  to  175020 => aso_source_data <= to_unsigned( 554 ,32);
when  175021  to  183269 => aso_source_data <= to_unsigned( 556 ,32);
when  183270  to  191906 => aso_source_data <= to_unsigned( 559 ,32);
when  191907  to  200950 => aso_source_data <= to_unsigned( 561 ,32);
when  200951  to  210421 => aso_source_data <= to_unsigned( 564 ,32);
when  210422  to  220338 => aso_source_data <= to_unsigned( 567 ,32);
when  220339  to  230722 => aso_source_data <= to_unsigned( 569 ,32);
when  230723  to  241596 => aso_source_data <= to_unsigned( 572 ,32);
when  241597  to  252982 => aso_source_data <= to_unsigned( 574 ,32);
when  252983  to  264904 => aso_source_data <= to_unsigned( 577 ,32);
when  264905  to  277389 => aso_source_data <= to_unsigned( 579 ,32);
when  277390  to  290462 => aso_source_data <= to_unsigned( 582 ,32);
when  290463  to  304151 => aso_source_data <= to_unsigned( 584 ,32);
when  304152  to  318485 => aso_source_data <= to_unsigned( 587 ,32);
when  318486  to  333495 => aso_source_data <= to_unsigned( 590 ,32);
when  333496  to  349212 => aso_source_data <= to_unsigned( 592 ,32);
when  349213  to  365670 => aso_source_data <= to_unsigned( 595 ,32);
when  365671  to  382904 => aso_source_data <= to_unsigned( 597 ,32);
when  382905  to  400949 => aso_source_data <= to_unsigned( 600 ,32);
when  400950  to  419845 => aso_source_data <= to_unsigned( 602 ,32);
when  419846  to  439632 => aso_source_data <= to_unsigned( 605 ,32);
when  439633  to  460351 => aso_source_data <= to_unsigned( 607 ,32);
when  460352  to  482047 => aso_source_data <= to_unsigned( 610 ,32);
when  482048  to  504765 => aso_source_data <= to_unsigned( 613 ,32);
when  504766  to  528554 => aso_source_data <= to_unsigned( 615 ,32);
when  528555  to  553464 => aso_source_data <= to_unsigned( 618 ,32);
when  553465  to  579548 => aso_source_data <= to_unsigned( 620 ,32);
when  579549  to  606862 => aso_source_data <= to_unsigned( 623 ,32);
when  606863  to  635462 => aso_source_data <= to_unsigned( 625 ,32);
when  635463  to  665411 => aso_source_data <= to_unsigned( 628 ,32);
when  665412  to  696770 => aso_source_data <= to_unsigned( 631 ,32);
when  696771  to  729608 => aso_source_data <= to_unsigned( 633 ,32);
when  729609  to  763994 => aso_source_data <= to_unsigned( 636 ,32);
when  763995  to  799999 => aso_source_data <= to_unsigned( 638 ,32);
when  800000  to  837702 => aso_source_data <= to_unsigned( 641 ,32);
when  837703  to  877182 => aso_source_data <= to_unsigned( 643 ,32);
when  877183  to  918522 => aso_source_data <= to_unsigned( 646 ,32);
when  918523  to  961811 => aso_source_data <= to_unsigned( 648 ,32);
when  961812  to  1007140 => aso_source_data <= to_unsigned( 651 ,32);
when  1007141  to  1054605 => aso_source_data <= to_unsigned( 654 ,32);
when  1054606  to  1104307 => aso_source_data <= to_unsigned( 656 ,32);
when  1104308  to  1156351 => aso_source_data <= to_unsigned( 659 ,32);
when  1156352  to  1210848 => aso_source_data <= to_unsigned( 661 ,32);
when  1210849  to  1267914 => aso_source_data <= to_unsigned( 664 ,32);
when  1267915  to  1327669 => aso_source_data <= to_unsigned( 666 ,32);
when  1327670  to  1390240 => aso_source_data <= to_unsigned( 669 ,32);
when  1390241  to  1455760 => aso_source_data <= to_unsigned( 671 ,32);
when  1455761  to  1524368 => aso_source_data <= to_unsigned( 674 ,32);
when  1524369  to  1596209 => aso_source_data <= to_unsigned( 677 ,32);
when  1596210  to  1671436 => aso_source_data <= to_unsigned( 679 ,32);
when  1671437  to  1750209 => aso_source_data <= to_unsigned( 682 ,32);
when  1750210  to  1832694 => aso_source_data <= to_unsigned( 684 ,32);
when  1832695  to  1919066 => aso_source_data <= to_unsigned( 687 ,32);
when  1919067  to  2009509 => aso_source_data <= to_unsigned( 689 ,32);
when  2009510  to  2104214 => aso_source_data <= to_unsigned( 692 ,32);
when  2104215  to  2203382 => aso_source_data <= to_unsigned( 695 ,32);
when  2203383  to  2307225 => aso_source_data <= to_unsigned( 697 ,32);
when  2307226  to  2415961 => aso_source_data <= to_unsigned( 700 ,32);
when  2415962  to  2529822 => aso_source_data <= to_unsigned( 702 ,32);
when  2529823  to  2649048 => aso_source_data <= to_unsigned( 705 ,32);
when  2649049  to  2773894 => aso_source_data <= to_unsigned( 707 ,32);
when  2773895  to  2904624 => aso_source_data <= to_unsigned( 710 ,32);
when  2904625  to  3041515 => aso_source_data <= to_unsigned( 712 ,32);
when  3041516  to  3184857 => aso_source_data <= to_unsigned( 715 ,32);
when  3184858  to  3334955 => aso_source_data <= to_unsigned( 718 ,32);
when  3334956  to  3492126 => aso_source_data <= to_unsigned( 720 ,32);
when  3492127  to  3656705 => aso_source_data <= to_unsigned( 723 ,32);
when  3656706  to  3829040 => aso_source_data <= to_unsigned( 725 ,32);
when  3829041  to  4009497 => aso_source_data <= to_unsigned( 728 ,32);
when  4009498  to  4198459 => aso_source_data <= to_unsigned( 730 ,32);
when  4198460  to  4396326 => aso_source_data <= to_unsigned( 733 ,32);
when  4396327  to  4603519 => aso_source_data <= to_unsigned( 735 ,32);
when  4603520  to  4820476 => aso_source_data <= to_unsigned( 738 ,32);
when  4820477  to  5047658 => aso_source_data <= to_unsigned( 741 ,32);
when  5047659  to  5285547 => aso_source_data <= to_unsigned( 743 ,32);
when  5285548  to  5534647 => aso_source_data <= to_unsigned( 746 ,32);
when  5534648  to  5795487 => aso_source_data <= to_unsigned( 748 ,32);
when  5795488  to  6068620 => aso_source_data <= to_unsigned( 751 ,32);
when  6068621  to  6354625 => aso_source_data <= to_unsigned( 753 ,32);
when  6354626  to  6654110 => aso_source_data <= to_unsigned( 756 ,32);
when  6654111  to  6967708 => aso_source_data <= to_unsigned( 759 ,32);
when  6967709  to  7296086 => aso_source_data <= to_unsigned( 761 ,32);
when  7296087  to  7639940 => aso_source_data <= to_unsigned( 764 ,32);
when  7639941  to  7999999 => aso_source_data <= to_unsigned( 766 ,32);
when  8000000  to  8377028 => aso_source_data <= to_unsigned( 769 ,32);
when  8377029  to  8771825 => aso_source_data <= to_unsigned( 771 ,32);
when  8771826  to  9185228 => aso_source_data <= to_unsigned( 774 ,32);
when  9185229  to  9618115 => aso_source_data <= to_unsigned( 776 ,32);
when  9618116  to  10071403 => aso_source_data <= to_unsigned( 779 ,32);
when  10071404  to  10546053 => aso_source_data <= to_unsigned( 782 ,32);
when  10546054  to  11043074 => aso_source_data <= to_unsigned( 784 ,32);
when  11043075  to  11563518 => aso_source_data <= to_unsigned( 787 ,32);
when  11563519  to  12108489 => aso_source_data <= to_unsigned( 789 ,32);
when  12108490  to  12679145 => aso_source_data <= to_unsigned( 792 ,32);
when  12679146  to  13276695 => aso_source_data <= to_unsigned( 794 ,32);
when  13276696  to  13902406 => aso_source_data <= to_unsigned( 797 ,32);
when  13902407  to  14557606 => aso_source_data <= to_unsigned( 799 ,32);
when  14557607  to  15243685 => aso_source_data <= to_unsigned( 802 ,32);
when  15243686  to  15962098 => aso_source_data <= to_unsigned( 805 ,32);
when  15962099  to  16714369 => aso_source_data <= to_unsigned( 807 ,32);
when  16714370  to  17502092 => aso_source_data <= to_unsigned( 810 ,32);
when  17502093  to  18326941 => aso_source_data <= to_unsigned( 812 ,32);
when  18326942  to  19190663 => aso_source_data <= to_unsigned( 815 ,32);
when  19190664  to  20095091 => aso_source_data <= to_unsigned( 817 ,32);
when  20095092  to  21042143 => aso_source_data <= to_unsigned( 820 ,32);
when  21042144  to  22033829 => aso_source_data <= to_unsigned( 823 ,32);
when  22033830  to  23072252 => aso_source_data <= to_unsigned( 825 ,32);
when  23072253  to  24159613 => aso_source_data <= to_unsigned( 828 ,32);
when  24159614  to  25298221 => aso_source_data <= to_unsigned( 830 ,32);
when  25298222  to  26490489 => aso_source_data <= to_unsigned( 833 ,32);
when  26490490  to  27738948 => aso_source_data <= to_unsigned( 835 ,32);
when  27738949  to  29046244 => aso_source_data <= to_unsigned( 838 ,32);
when  29046245  to  30415151 => aso_source_data <= to_unsigned( 840 ,32);
when  30415152  to  31848573 => aso_source_data <= to_unsigned( 843 ,32);
when  31848574  to  33349550 => aso_source_data <= to_unsigned( 846 ,32);
when  33349551  to  34921266 => aso_source_data <= to_unsigned( 848 ,32);
when  34921267  to  36567055 => aso_source_data <= to_unsigned( 851 ,32);
when  36567056  to  38290407 => aso_source_data <= to_unsigned( 853 ,32);
when  38290408  to  40094978 => aso_source_data <= to_unsigned( 856 ,32);
when  40094979  to  41984596 => aso_source_data <= to_unsigned( 858 ,32);
when  41984597  to  43963269 => aso_source_data <= to_unsigned( 861 ,32);
when  43963270  to  46035194 => aso_source_data <= to_unsigned( 863 ,32);
when  46035195  to  48204766 => aso_source_data <= to_unsigned( 866 ,32);
when  48204767  to  50476587 => aso_source_data <= to_unsigned( 869 ,32);
when  50476588  to  52855475 => aso_source_data <= to_unsigned( 871 ,32);
when  52855476  to  55346477 => aso_source_data <= to_unsigned( 874 ,32);
when  55346478  to  57954876 => aso_source_data <= to_unsigned( 876 ,32);
when  57954877  to  60686206 => aso_source_data <= to_unsigned( 879 ,32);
when  60686207  to  63546258 => aso_source_data <= to_unsigned( 881 ,32);
when  63546259  to  66541101 => aso_source_data <= to_unsigned( 884 ,32);
when  66541102  to  69677087 => aso_source_data <= to_unsigned( 887 ,32);
when  69677088  to  72960867 => aso_source_data <= to_unsigned( 889 ,32);
when  72960868  to  76399406 => aso_source_data <= to_unsigned( 892 ,32);
when  76399407  to  79999999 => aso_source_data <= to_unsigned( 894 ,32);
when  80000000  to  83770283 => aso_source_data <= to_unsigned( 897 ,32);
when  83770284  to  87718255 => aso_source_data <= to_unsigned( 899 ,32);
when  87718256  to  91852289 => aso_source_data <= to_unsigned( 902 ,32);
when  91852290  to  96181154 => aso_source_data <= to_unsigned( 904 ,32);
when  96181155  to  100714032 => aso_source_data <= to_unsigned( 907 ,32);
when  100714033  to  105460539 => aso_source_data <= to_unsigned( 910 ,32);
when  105460540  to  110430741 => aso_source_data <= to_unsigned( 912 ,32);
when  110430742  to  115635181 => aso_source_data <= to_unsigned( 915 ,32);
when  115635182  to  121084899 => aso_source_data <= to_unsigned( 917 ,32);
when  121084900  to  126791455 => aso_source_data <= to_unsigned( 920 ,32);
when  126791456  to  132766952 => aso_source_data <= to_unsigned( 922 ,32);
when  132766953  to  139024066 => aso_source_data <= to_unsigned( 925 ,32);
when  139024067  to  145576068 => aso_source_data <= to_unsigned( 927 ,32);
when  145576069  to  152436857 => aso_source_data <= to_unsigned( 930 ,32);
when  152436858  to  159620985 => aso_source_data <= to_unsigned( 933 ,32);
when  159620986  to  167143690 => aso_source_data <= to_unsigned( 935 ,32);
when  167143691  to  175020929 => aso_source_data <= to_unsigned( 938 ,32);
when  175020930  to  183269412 => aso_source_data <= to_unsigned( 940 ,32);
when  183269413  to  191906633 => aso_source_data <= to_unsigned( 943 ,32);
when  191906634  to  200950914 => aso_source_data <= to_unsigned( 945 ,32);
when  200950915  to  210421439 => aso_source_data <= to_unsigned( 948 ,32);
when  210421440  to  220338296 => aso_source_data <= to_unsigned( 951 ,32);
when  220338297  to  230722520 => aso_source_data <= to_unsigned( 953 ,32);
when  230722521  to  241596137 => aso_source_data <= to_unsigned( 956 ,32);
when  241596138  to  252982212 => aso_source_data <= to_unsigned( 958 ,32);
when  252982213  to  264904897 => aso_source_data <= to_unsigned( 961 ,32);
when  264904898  to  277389480 => aso_source_data <= to_unsigned( 963 ,32);
when  277389481  to  290462443 => aso_source_data <= to_unsigned( 966 ,32);
when  290462444  to  304151517 => aso_source_data <= to_unsigned( 968 ,32);
when  304151518  to  318485736 => aso_source_data <= to_unsigned( 971 ,32);
when  318485737  to  333495506 => aso_source_data <= to_unsigned( 974 ,32);
when  333495507  to  349212665 => aso_source_data <= to_unsigned( 976 ,32);
when  349212666  to  365670551 => aso_source_data <= to_unsigned( 979 ,32);
when  365670552  to  382904073 => aso_source_data <= to_unsigned( 981 ,32);
when  382904074  to  400949786 => aso_source_data <= to_unsigned( 984 ,32);
when  400949787  to  419845968 => aso_source_data <= to_unsigned( 986 ,32);
when  419845969  to  439632699 => aso_source_data <= to_unsigned( 989 ,32);
when  439632700  to  460351949 => aso_source_data <= to_unsigned( 991 ,32);
when  460351950  to  482047668 => aso_source_data <= to_unsigned( 994 ,32);
when  482047669  to  504765875 => aso_source_data <= to_unsigned( 997 ,32);
when  504765876  to  528554758 => aso_source_data <= to_unsigned( 999 ,32);
when  528554759  to  553464776 => aso_source_data <= to_unsigned( 1002 ,32);
when  553464777  to  579548768 => aso_source_data <= to_unsigned( 1004 ,32);
when  579548769  to  606862060 => aso_source_data <= to_unsigned( 1007 ,32);
when  606862061  to  635462587 => aso_source_data <= to_unsigned( 1009 ,32);
when  635462588  to  665411016 => aso_source_data <= to_unsigned( 1012 ,32);
when  665411017  to  696770871 => aso_source_data <= to_unsigned( 1015 ,32);
when  696770872  to  729608671 => aso_source_data <= to_unsigned( 1017 ,32);
when  729608672  to  763994068 => aso_source_data <= to_unsigned( 1020 ,32);
when  763994069  to  799999999 => aso_source_data <= to_unsigned( 1022 ,32);
when  800000000  to  837702838 => aso_source_data <= to_unsigned( 1025 ,32);
when  837702839  to  877182556 => aso_source_data <= to_unsigned( 1027 ,32);
when  877182557  to  918522897 => aso_source_data <= to_unsigned( 1030 ,32);
when  918522898  to  961811547 => aso_source_data <= to_unsigned( 1032 ,32);
when  961811548  to  1007140329 => aso_source_data <= to_unsigned( 1035 ,32);
when  1007140330  to  1054605390 => aso_source_data <= to_unsigned( 1038 ,32);
when  1054605391  to  1104307411 => aso_source_data <= to_unsigned( 1040 ,32);
when  1104307412  to  1156351816 => aso_source_data <= to_unsigned( 1043 ,32);
when  1156351817  to  1210848998 => aso_source_data <= to_unsigned( 1045 ,32);
when  1210848999  to  1267914553 => aso_source_data <= to_unsigned( 1048 ,32);
when  1267914554  to  1327669525 => aso_source_data <= to_unsigned( 1050 ,32);
when  1327669526  to  1390240662 => aso_source_data <= to_unsigned( 1053 ,32);
when  1390240663  to  1455760686 => aso_source_data <= to_unsigned( 1055 ,32);
when  1455760687  to  1524368574 => aso_source_data <= to_unsigned( 1058 ,32);
when  1524368575  to  1596209851 => aso_source_data <= to_unsigned( 1061 ,32);
when  1596209852  to  1671436904 => aso_source_data <= to_unsigned( 1063 ,32);
when  1671436905  to  1750209299 => aso_source_data <= to_unsigned( 1066 ,32);
when  1750209300  to  1832694122 => aso_source_data <= to_unsigned( 1068 ,32);
when  1832694123  to  1919066335 => aso_source_data <= to_unsigned( 1071 ,32);
when  1919066336  to  2009509145 => aso_source_data <= to_unsigned( 1073 ,32);
when  2009509146  to  2104214393 => aso_source_data <= to_unsigned( 1076 ,32);
when others => aso_source_data <= (others => '0');
			
			end case;
		end if;
    end process;
o_bit_index <= bit_fft_index;
end behav;